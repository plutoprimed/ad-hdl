//
// generated from this migen source: https://github.com/m-labs/cossin/blob/master/cossin.ipynb
//

/* Machine-generated using Migen */
module cossin(
	input [17:0] z,
	output signed [15:0] x,
	output signed [15:0] y,
	input clk
);

wire [14:0] lut_x;
wire [14:0] lut_y;
wire [2:0] lut_xd;
wire [2:0] lut_yd;
wire [8:0] adr;
wire [35:0] dat_r;
wire [14:0] za;
wire signed [5:0] zd;
wire signed [5:0] zd_cossingen0;
reg signed [5:0] zd_cossingen1 = 6'sd0;
reg signed [5:0] zd_cossingen2 = 6'sd0;
wire [2:0] zq_cossingen0;
reg [2:0] zq_cossingen1 = 3'd0;
reg [2:0] zq_cossingen2 = 3'd0;
wire signed [15:0] x1;
wire signed [15:0] y1;
wire signed [15:0] x2;
wire signed [15:0] y2;
wire [35:0] cossingen0;
reg [35:0] cossingen1 = 36'd0;

// synthesis translate_off
reg dummy_s;
initial dummy_s <= 1'd0;
// synthesis translate_on

assign zd = (za[5:0] - 6'd32);
assign zd_cossingen0 = zd;
assign zq_cossingen0 = {z[17], (z[16] ^ z[17]), (z[15] ^ z[16])};
assign cossingen0 = dat_r;
assign za = (z[15] ? (15'd32767 - z[14:0]) : z[14:0]);
assign adr = za[14:6];
assign {lut_yd, lut_xd, lut_y, lut_x} = cossingen1;
assign x1 = ($signed({1'd0, lut_x}) - (((zd_cossingen2 * $signed({1'd0, lut_yd})) + $signed({1'd0, 3'd4})) >>> 2'd3));
assign y1 = ($signed({1'd0, lut_y}) + (((zd_cossingen2 * $signed({1'd0, lut_xd})) + $signed({1'd0, 3'd4})) >>> 2'd3));
assign x2 = (zq_cossingen2[0] ? y1 : x1);
assign y2 = (zq_cossingen2[0] ? x1 : y1);
assign x = (zq_cossingen2[1] ? (-x2) : x2);
assign y = (zq_cossingen2[2] ? (-y2) : y2);

always @(posedge clk) begin
	zd_cossingen1 <= zd_cossingen0;
	zd_cossingen2 <= zd_cossingen1;
	zq_cossingen1 <= zq_cossingen0;
	zq_cossingen2 <= zq_cossingen1;
	cossingen1 <= cossingen0;
end

reg [35:0] mem[0:511];
reg [8:0] memadr;
always @(posedge clk) begin
	memadr <= adr;
end

assign dat_r = mem[memadr];

initial begin
    mem [0] = 36'h1800cffff;
    mem [1] = 36'h18025ffff;
    mem [2] = 36'h1803f7fff;
    mem [3] = 36'h180587fff;
    mem [4] = 36'h180717ffe;
    mem [5] = 36'h1808a7ffe;
    mem [6] = 36'h180a3fffd;
    mem [7] = 36'h180bcfffd;
    mem [8] = 36'h180d5fffc;
    mem [9] = 36'h180eefffc;
    mem [10] = 36'h181087ffb;
    mem [11] = 36'h181217ffa;
    mem [12] = 36'h1813a7ff9;
    mem [13] = 36'h18153fff8;
    mem [14] = 36'h1816cfff7;
    mem [15] = 36'h18185fff6;
    mem [16] = 36'h1819efff5;
    mem [17] = 36'h181b87ff3;
    mem [18] = 36'h181d17ff2;
    mem [19] = 36'h181ea7ff0;
    mem [20] = 36'h182037fef;
    mem [21] = 36'h1821c7fed;
    mem [22] = 36'h18235ffeb;
    mem [23] = 36'h1824effea;
    mem [24] = 36'h18267ffe8;
    mem [25] = 36'h18280ffe6;
    mem [26] = 36'h1829a7fe4;
    mem [27] = 36'h182b37fe2;
    mem [28] = 36'h182cc7fe0;
    mem [29] = 36'h182e57fdd;
    mem [30] = 36'h182fe7fdb;
    mem [31] = 36'h18317ffd9;
    mem [32] = 36'h18330ffd6;
    mem [33] = 36'h18349ffd4;
    mem [34] = 36'h18362ffd1;
    mem [35] = 36'h1837bffce;
    mem [36] = 36'h183957fcc;
    mem [37] = 36'h183ae7fc9;
    mem [38] = 36'h183c77fc6;
    mem [39] = 36'h183e07fc3;
    mem [40] = 36'h183f97fc0;
    mem [41] = 36'h18412ffbd;
    mem [42] = 36'h1842bffb9;
    mem [43] = 36'h18444ffb6;
    mem [44] = 36'h1845dffb3;
    mem [45] = 36'h18476ffaf;
    mem [46] = 36'h1848fffac;
    mem [47] = 36'h184a8ffa8;
    mem [48] = 36'h184c27fa4;
    mem [49] = 36'h184db7fa1;
    mem [50] = 36'h184f47f9d;
    mem [51] = 36'h1850d7f99;
    mem [52] = 36'h385267f95;
    mem [53] = 36'h3853f7f91;
    mem [54] = 36'h385587f8d;
    mem [55] = 36'h385717f88;
    mem [56] = 36'h3858a7f84;
    mem [57] = 36'h385a37f80;
    mem [58] = 36'h385bc7f7b;
    mem [59] = 36'h385d5ff77;
    mem [60] = 36'h385eeff72;
    mem [61] = 36'h38607ff6d;
    mem [62] = 36'h38620ff69;
    mem [63] = 36'h38639ff64;
    mem [64] = 36'h38652ff5f;
    mem [65] = 36'h3866bff5a;
    mem [66] = 36'h38684ff55;
    mem [67] = 36'h3869dff50;
    mem [68] = 36'h386b6ff4a;
    mem [69] = 36'h386cfff45;
    mem [70] = 36'h386e8ff40;
    mem [71] = 36'h38701ff3a;
    mem [72] = 36'h3871aff35;
    mem [73] = 36'h38733ff2f;
    mem [74] = 36'h3874cff29;
    mem [75] = 36'h387657f23;
    mem [76] = 36'h3877e7f1e;
    mem [77] = 36'h387977f18;
    mem [78] = 36'h387b07f12;
    mem [79] = 36'h387c97f0c;
    mem [80] = 36'h387e27f05;
    mem [81] = 36'h387fb7eff;
    mem [82] = 36'h388147ef9;
    mem [83] = 36'h3882d7ef3;
    mem [84] = 36'h38845feec;
    mem [85] = 36'h3885efee6;
    mem [86] = 36'h38877fedf;
    mem [87] = 36'h38890fed8;
    mem [88] = 36'h388a9fed2;
    mem [89] = 36'h388c2fecb;
    mem [90] = 36'h388db7ec4;
    mem [91] = 36'h388f47ebd;
    mem [92] = 36'h3890d7eb6;
    mem [93] = 36'h389267eaf;
    mem [94] = 36'h3893efea7;
    mem [95] = 36'h38957fea0;
    mem [96] = 36'h38970fe99;
    mem [97] = 36'h389897e91;
    mem [98] = 36'h389a27e8a;
    mem [99] = 36'h389bb7e82;
    mem [100] = 36'h389d47e7a;
    mem [101] = 36'h389ecfe73;
    mem [102] = 36'h38a05fe6b;
    mem [103] = 36'h38a1e7e63;
    mem [104] = 36'h38a377e5b;
    mem [105] = 36'h38a507e53;
    mem [106] = 36'h38a68fe4b;
    mem [107] = 36'h38a81fe42;
    mem [108] = 36'h38a9a7e3a;
    mem [109] = 36'h38ab37e32;
    mem [110] = 36'h38acc7e29;
    mem [111] = 36'h38ae4fe21;
    mem [112] = 36'h38afdfe18;
    mem [113] = 36'h38b167e10;
    mem [114] = 36'h38b2f7e07;
    mem [115] = 36'h38b47fdfe;
    mem [116] = 36'h38b60fdf5;
    mem [117] = 36'h38b797dec;
    mem [118] = 36'h38b927de3;
    mem [119] = 36'h38baafdda;
    mem [120] = 36'h38bc37dd1;
    mem [121] = 36'h38bdc7dc8;
    mem [122] = 36'h38bf4fdbe;
    mem [123] = 36'h38c0dfdb5;
    mem [124] = 36'h38c267dab;
    mem [125] = 36'h38c3efda2;
    mem [126] = 36'h38c57fd98;
    mem [127] = 36'h38c707d8e;
    mem [128] = 36'h38c88fd84;
    mem [129] = 36'h38ca17d7b;
    mem [130] = 36'h38cba7d71;
    mem [131] = 36'h38cd2fd67;
    mem [132] = 36'h38ceb7d5c;
    mem [133] = 36'h38d03fd52;
    mem [134] = 36'h38d1cfd48;
    mem [135] = 36'h38d357d3e;
    mem [136] = 36'h38d4dfd33;
    mem [137] = 36'h38d667d29;
    mem [138] = 36'h38d7efd1e;
    mem [139] = 36'h38d977d14;
    mem [140] = 36'h38db07d09;
    mem [141] = 36'h38dc8fcfe;
    mem [142] = 36'h38de17cf3;
    mem [143] = 36'h38df9fce8;
    mem [144] = 36'h38e127cdd;
    mem [145] = 36'h38e2afcd2;
    mem [146] = 36'h38e437cc7;
    mem [147] = 36'h38e5bfcbc;
    mem [148] = 36'h38e747cb1;
    mem [149] = 36'h38e8cfca5;
    mem [150] = 36'h38ea57c9a;
    mem [151] = 36'h38ebdfc8e;
    mem [152] = 36'h38ed67c83;
    mem [153] = 36'h38eee7c77;
    mem [154] = 36'h38f06fc6b;
    mem [155] = 36'h38f1f7c5f;
    mem [156] = 36'h38f37fc53;
    mem [157] = 36'h58f507c47;
    mem [158] = 36'h58f68fc3b;
    mem [159] = 36'h58f80fc2f;
    mem [160] = 36'h58f997c23;
    mem [161] = 36'h58fb1fc17;
    mem [162] = 36'h58fca7c0a;
    mem [163] = 36'h58fe27bfe;
    mem [164] = 36'h58ffafbf1;
    mem [165] = 36'h590137be5;
    mem [166] = 36'h5902b7bd8;
    mem [167] = 36'h59043fbcb;
    mem [168] = 36'h5905bfbbf;
    mem [169] = 36'h590747bb2;
    mem [170] = 36'h5908cfba5;
    mem [171] = 36'h590a4fb98;
    mem [172] = 36'h590bd7b8b;
    mem [173] = 36'h590d57b7d;
    mem [174] = 36'h590edfb70;
    mem [175] = 36'h59105fb63;
    mem [176] = 36'h5911e7b55;
    mem [177] = 36'h591367b48;
    mem [178] = 36'h5914e7b3a;
    mem [179] = 36'h59166fb2d;
    mem [180] = 36'h5917efb1f;
    mem [181] = 36'h591977b11;
    mem [182] = 36'h591af7b03;
    mem [183] = 36'h591c77af5;
    mem [184] = 36'h591df7ae7;
    mem [185] = 36'h591f7fad9;
    mem [186] = 36'h5920ffacb;
    mem [187] = 36'h59227fabd;
    mem [188] = 36'h5923ffaaf;
    mem [189] = 36'h59257faa0;
    mem [190] = 36'h592707a92;
    mem [191] = 36'h592887a83;
    mem [192] = 36'h592a07a75;
    mem [193] = 36'h592b87a66;
    mem [194] = 36'h592d07a57;
    mem [195] = 36'h592e87a49;
    mem [196] = 36'h593007a3a;
    mem [197] = 36'h593187a2b;
    mem [198] = 36'h593307a1c;
    mem [199] = 36'h593487a0d;
    mem [200] = 36'h5936079fd;
    mem [201] = 36'h5937879ee;
    mem [202] = 36'h5939079df;
    mem [203] = 36'h593a7f9cf;
    mem [204] = 36'h593bff9c0;
    mem [205] = 36'h593d7f9b0;
    mem [206] = 36'h593eff9a1;
    mem [207] = 36'h59407f991;
    mem [208] = 36'h5941f7981;
    mem [209] = 36'h594377971;
    mem [210] = 36'h5944f7962;
    mem [211] = 36'h59466f952;
    mem [212] = 36'h5947ef941;
    mem [213] = 36'h59496f931;
    mem [214] = 36'h594ae7921;
    mem [215] = 36'h594c67911;
    mem [216] = 36'h594ddf901;
    mem [217] = 36'h594f5f8f0;
    mem [218] = 36'h5950d78e0;
    mem [219] = 36'h5952578cf;
    mem [220] = 36'h5953cf8be;
    mem [221] = 36'h5955478ae;
    mem [222] = 36'h5956c789d;
    mem [223] = 36'h59583f88c;
    mem [224] = 36'h5959bf87b;
    mem [225] = 36'h595b3786a;
    mem [226] = 36'h595caf859;
    mem [227] = 36'h595e27848;
    mem [228] = 36'h595fa7837;
    mem [229] = 36'h59611f825;
    mem [230] = 36'h596297814;
    mem [231] = 36'h59640f803;
    mem [232] = 36'h5965877f1;
    mem [233] = 36'h5966ff7df;
    mem [234] = 36'h5968777ce;
    mem [235] = 36'h5969ef7bc;
    mem [236] = 36'h596b677aa;
    mem [237] = 36'h596cdf798;
    mem [238] = 36'h596e57786;
    mem [239] = 36'h596fcf774;
    mem [240] = 36'h597147762;
    mem [241] = 36'h5972bf750;
    mem [242] = 36'h59743773e;
    mem [243] = 36'h5975af72c;
    mem [244] = 36'h59771f719;
    mem [245] = 36'h597897707;
    mem [246] = 36'h597a0f6f4;
    mem [247] = 36'h597b876e2;
    mem [248] = 36'h597cf76cf;
    mem [249] = 36'h597e6f6bc;
    mem [250] = 36'h597fe76a9;
    mem [251] = 36'h598157697;
    mem [252] = 36'h5982cf684;
    mem [253] = 36'h59843f671;
    mem [254] = 36'h5985b765e;
    mem [255] = 36'h59872764a;
    mem [256] = 36'h59889f637;
    mem [257] = 36'h598a0f624;
    mem [258] = 36'h598b7f610;
    mem [259] = 36'h598cf75fd;
    mem [260] = 36'h598e675e9;
    mem [261] = 36'h598fd75d6;
    mem [262] = 36'h59914f5c2;
    mem [263] = 36'h5992bf5ae;
    mem [264] = 36'h59942f59b;
    mem [265] = 36'h59959f587;
    mem [266] = 36'h59970f573;
    mem [267] = 36'h79987f55f;
    mem [268] = 36'h7999f754b;
    mem [269] = 36'h799b67537;
    mem [270] = 36'h799cd7522;
    mem [271] = 36'h799e4750e;
    mem [272] = 36'h799fb74fa;
    mem [273] = 36'h79a11f4e5;
    mem [274] = 36'h79a28f4d1;
    mem [275] = 36'h79a3ff4bc;
    mem [276] = 36'h79a56f4a8;
    mem [277] = 36'h79a6df493;
    mem [278] = 36'h79a84f47e;
    mem [279] = 36'h79a9b7469;
    mem [280] = 36'h79ab27454;
    mem [281] = 36'h79ac9743f;
    mem [282] = 36'h79adff42a;
    mem [283] = 36'h79af6f415;
    mem [284] = 36'h79b0d7400;
    mem [285] = 36'h79b2473eb;
    mem [286] = 36'h79b3b73d5;
    mem [287] = 36'h79b51f3c0;
    mem [288] = 36'h79b6873aa;
    mem [289] = 36'h79b7f7395;
    mem [290] = 36'h79b95f37f;
    mem [291] = 36'h79bacf369;
    mem [292] = 36'h79bc37354;
    mem [293] = 36'h79bd9f33e;
    mem [294] = 36'h79bf07328;
    mem [295] = 36'h79c077312;
    mem [296] = 36'h79c1df2fc;
    mem [297] = 36'h79c3472e6;
    mem [298] = 36'h79c4af2d0;
    mem [299] = 36'h79c6172b9;
    mem [300] = 36'h79c77f2a3;
    mem [301] = 36'h79c8e728d;
    mem [302] = 36'h79ca4f276;
    mem [303] = 36'h79cbb7260;
    mem [304] = 36'h79cd1f249;
    mem [305] = 36'h79ce87232;
    mem [306] = 36'h79cfef21c;
    mem [307] = 36'h79d14f205;
    mem [308] = 36'h79d2b71ee;
    mem [309] = 36'h79d41f1d7;
    mem [310] = 36'h79d5871c0;
    mem [311] = 36'h79d6e71a9;
    mem [312] = 36'h79d84f192;
    mem [313] = 36'h79d9af17a;
    mem [314] = 36'h79db17163;
    mem [315] = 36'h79dc7714c;
    mem [316] = 36'h79dddf134;
    mem [317] = 36'h79df3f11d;
    mem [318] = 36'h79e0a7105;
    mem [319] = 36'h79e2070ee;
    mem [320] = 36'h79e3670d6;
    mem [321] = 36'h79e4cf0be;
    mem [322] = 36'h79e62f0a6;
    mem [323] = 36'h79e78f08f;
    mem [324] = 36'h79e8ef077;
    mem [325] = 36'h79ea5705f;
    mem [326] = 36'h79ebb7046;
    mem [327] = 36'h79ed1702e;
    mem [328] = 36'h79ee77016;
    mem [329] = 36'h75efd6ffe;
    mem [330] = 36'h75f136fe5;
    mem [331] = 36'h75f296fcd;
    mem [332] = 36'h75f3eefb4;
    mem [333] = 36'h75f54ef9c;
    mem [334] = 36'h75f6aef83;
    mem [335] = 36'h75f80ef6b;
    mem [336] = 36'h75f96ef52;
    mem [337] = 36'h75fac6f39;
    mem [338] = 36'h75fc26f20;
    mem [339] = 36'h75fd86f07;
    mem [340] = 36'h75fedeeee;
    mem [341] = 36'h76003eed5;
    mem [342] = 36'h760196ebc;
    mem [343] = 36'h7602f6ea2;
    mem [344] = 36'h76044ee89;
    mem [345] = 36'h7605aee70;
    mem [346] = 36'h760706e56;
    mem [347] = 36'h76085ee3d;
    mem [348] = 36'h7609b6e23;
    mem [349] = 36'h760b16e0a;
    mem [350] = 36'h760c6edf0;
    mem [351] = 36'h760dc6dd6;
    mem [352] = 36'h760f1edbc;
    mem [353] = 36'h761076da2;
    mem [354] = 36'h7611ced88;
    mem [355] = 36'h761326d6e;
    mem [356] = 36'h76147ed54;
    mem [357] = 36'h7615d6d3a;
    mem [358] = 36'h76172ed20;
    mem [359] = 36'h761886d06;
    mem [360] = 36'h7619deceb;
    mem [361] = 36'h761b2ecd1;
    mem [362] = 36'h761c86cb6;
    mem [363] = 36'h761ddec9c;
    mem [364] = 36'h761f2ec81;
    mem [365] = 36'h762086c66;
    mem [366] = 36'h7621dec4c;
    mem [367] = 36'h76232ec31;
    mem [368] = 36'h76247ec16;
    mem [369] = 36'h7625d6bfb;
    mem [370] = 36'h762726be0;
    mem [371] = 36'h76287ebc5;
    mem [372] = 36'h7629cebaa;
    mem [373] = 36'h762b1eb8e;
    mem [374] = 36'h762c6eb73;
    mem [375] = 36'h762dc6b58;
    mem [376] = 36'h762f16b3c;
    mem [377] = 36'h763066b21;
    mem [378] = 36'h7631b6b05;
    mem [379] = 36'h763306aea;
    mem [380] = 36'h763456ace;
    mem [381] = 36'h7635a6ab2;
    mem [382] = 36'h7636f6a97;
    mem [383] = 36'h76383ea7b;
    mem [384] = 36'h76398ea5f;
    mem [385] = 36'h963adea43;
    mem [386] = 36'h963c2ea27;
    mem [387] = 36'h963d76a0b;
    mem [388] = 36'h963ec69ee;
    mem [389] = 36'h9640169d2;
    mem [390] = 36'h96415e9b6;
    mem [391] = 36'h9642ae99a;
    mem [392] = 36'h9643f697d;
    mem [393] = 36'h96453e961;
    mem [394] = 36'h96468e944;
    mem [395] = 36'h9647d6927;
    mem [396] = 36'h96491e90b;
    mem [397] = 36'h964a6e8ee;
    mem [398] = 36'h964bb68d1;
    mem [399] = 36'h964cfe8b4;
    mem [400] = 36'h964e46897;
    mem [401] = 36'h964f8e87a;
    mem [402] = 36'h9650d685d;
    mem [403] = 36'h96521e840;
    mem [404] = 36'h965366823;
    mem [405] = 36'h9654ae806;
    mem [406] = 36'h9655f67e8;
    mem [407] = 36'h9657367cb;
    mem [408] = 36'h96587e7ae;
    mem [409] = 36'h9659c6790;
    mem [410] = 36'h965b0e772;
    mem [411] = 36'h965c4e755;
    mem [412] = 36'h965d96737;
    mem [413] = 36'h965ed6719;
    mem [414] = 36'h96601e6fc;
    mem [415] = 36'h96615e6de;
    mem [416] = 36'h96629e6c0;
    mem [417] = 36'h9663e66a2;
    mem [418] = 36'h966526684;
    mem [419] = 36'h966666666;
    mem [420] = 36'h9667a6647;
    mem [421] = 36'h9668ee629;
    mem [422] = 36'h966a2e60b;
    mem [423] = 36'h966b6e5ec;
    mem [424] = 36'h966cae5ce;
    mem [425] = 36'h966dee5af;
    mem [426] = 36'h966f2e591;
    mem [427] = 36'h96706e572;
    mem [428] = 36'h9671a6554;
    mem [429] = 36'h9672e6535;
    mem [430] = 36'h967426516;
    mem [431] = 36'h96755e4f7;
    mem [432] = 36'h96769e4d8;
    mem [433] = 36'h9677de4b9;
    mem [434] = 36'h96791649a;
    mem [435] = 36'h967a5647b;
    mem [436] = 36'h967b8e45c;
    mem [437] = 36'h967cce43d;
    mem [438] = 36'h967e0641d;
    mem [439] = 36'h967f3e3fe;
    mem [440] = 36'h9680763df;
    mem [441] = 36'h9681b63bf;
    mem [442] = 36'h9682ee3a0;
    mem [443] = 36'h968426380;
    mem [444] = 36'h96855e360;
    mem [445] = 36'h968696341;
    mem [446] = 36'h9687ce321;
    mem [447] = 36'h968906301;
    mem [448] = 36'h968a3e2e1;
    mem [449] = 36'h968b6e2c1;
    mem [450] = 36'h968ca62a1;
    mem [451] = 36'h968dde281;
    mem [452] = 36'h968f16261;
    mem [453] = 36'h969046241;
    mem [454] = 36'h96917e221;
    mem [455] = 36'h9692ae200;
    mem [456] = 36'h9693e61e0;
    mem [457] = 36'h9695161c0;
    mem [458] = 36'h96964619f;
    mem [459] = 36'h96977e17f;
    mem [460] = 36'h9698ae15e;
    mem [461] = 36'h9699de13d;
    mem [462] = 36'h969b0e11d;
    mem [463] = 36'h969c3e0fc;
    mem [464] = 36'h969d760db;
    mem [465] = 36'h969ea60ba;
    mem [466] = 36'h969fd6099;
    mem [467] = 36'h96a0fe078;
    mem [468] = 36'h96a22e057;
    mem [469] = 36'h96a35e036;
    mem [470] = 36'h96a48e015;
    mem [471] = 36'h96a5bdff4;
    mem [472] = 36'h96a6e5fd2;
    mem [473] = 36'h96a815fb1;
    mem [474] = 36'h96a93df90;
    mem [475] = 36'h96aa6df6e;
    mem [476] = 36'h96ab95f4d;
    mem [477] = 36'h96acc5f2b;
    mem [478] = 36'h96adedf09;
    mem [479] = 36'h96af15ee8;
    mem [480] = 36'h96b045ec6;
    mem [481] = 36'h96b16dea4;
    mem [482] = 36'h96b295e82;
    mem [483] = 36'h96b3bde60;
    mem [484] = 36'h96b4e5e3e;
    mem [485] = 36'h96b60de1c;
    mem [486] = 36'h96b735dfa;
    mem [487] = 36'h96b85ddd8;
    mem [488] = 36'h96b985db6;
    mem [489] = 36'h96baa5d94;
    mem [490] = 36'h96bbcdd71;
    mem [491] = 36'h96bcf5d4f;
    mem [492] = 36'h96be15d2c;
    mem [493] = 36'h96bf3dd0a;
    mem [494] = 36'h96c065ce7;
    mem [495] = 36'h96c185cc5;
    mem [496] = 36'h96c2a5ca2;
    mem [497] = 36'h96c3cdc7f;
    mem [498] = 36'h96c4edc5d;
    mem [499] = 36'h96c60dc3a;
    mem [500] = 36'h96c72dc17;
    mem [501] = 36'h96c855bf4;
    mem [502] = 36'h96c975bd1;
    mem [503] = 36'h96ca95bae;
    mem [504] = 36'h92cbb5b8b;
    mem [505] = 36'h92ccd5b68;
    mem [506] = 36'h92cdedb44;
    mem [507] = 36'h92cf0db21;
    mem [508] = 36'h92d02dafe;
    mem [509] = 36'h92d14dada;
    mem [510] = 36'h92d265ab7;
    mem [511] = 36'h92d385a94;
end

endmodule

